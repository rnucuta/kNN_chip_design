parameter CLK_PERIOD = 440;        // Change based on timing violations from sdf backannotation
parameter PIPE_STAGES = 7;       // Change based on how long it takes to get first output
parameter DSIZE = 12; 			// bit size of dist accumulation (the sum of subdists)
